module isNotEqual_gate32(out, x, y);
	output out;
	input [31:0] x,y;
	wire [31:0] a;
	wire [15:0] b;
	wire [7:0] c;
	wire [3:0] d;
	wire [1:0] e;
	
	
	xor n0(a[0], x[0], y[0]);
	xor n1(a[1], x[1],y[1]);
	xor n2(a[2], x[2],y[2]);
	xor n3(a[3], x[3],y[3]);
	xor n4(a[4], x[4],y[4]);
	xor n5(a[5], x[5],y[5]);
	xor n6(a[6], x[6],y[6]);
	xor n7(a[7], x[7],y[7]);
	xor n8(a[8], x[8],y[8]);
	xor n9(a[9], x[9],y[9]);
	xor n10(a[10], x[10],y[10]);
	xor n11(a[11], x[11],y[11]);
	xor n12(a[12], x[12],y[12]);
	xor n13(a[13], x[13],y[13]);
	xor n14(a[14], x[14],y[14]);
	xor n15(a[15], x[15],y[15]);
	
	xor n16(a[16], x[16],y[16]);
	xor n17(a[17], x[17],y[17]);
	xor n18(a[18], x[18],y[18]);
	xor n19(a[19], x[19],y[19]);
	xor n20(a[20], x[20],y[20]);
	xor n21(a[21], x[21],y[21]);
	xor n22(a[22], x[22],y[22]);
	xor n23(a[23], x[23],y[23]);
	xor n24(a[24], x[24],y[24]);
	xor n25(a[25], x[25],y[25]);
	xor n26(a[26], x[26],y[26]);
	xor n27(a[27], x[27],y[27]);
	xor n28(a[28], x[28],y[28]);
	xor n29(a[29], x[29],y[29]);
	xor n30(a[30], x[30],y[30]);
	xor n31(a[31], x[31],y[31]);
	
	or n00(b[0], a[0], a[1]);
	or n01(b[1], a[3],a[2]);
	or n02(b[2], a[4],a[5]);
	or n03(b[3], a[6],a[7]);
	or n04(b[4], a[8],a[9]);
	or n05(b[5], a[10],a[11]);
	or n06(b[6], a[12],a[13]);
	or n07(b[7], a[14],a[15]);
	or n08(b[8], a[16],a[17]);
	or n09(b[9], a[18],a[19]);
	or n010(b[10], a[20],a[21]);
	or n011(b[11], a[22],a[23]);
	or n012(b[12], a[24],a[25]);
	or n013(b[13], a[26],a[27]);
	or n014(b[14], a[28],a[29]);
	or n015(b[15], a[30],a[31]);
	
	or n000(c[0], b[0], b[1]);
	or n001(c[1], b[3], b[2]);
	or n002(c[2], b[4], b[5]);
	or n003(c[3], b[6], b[7]);
	or n004(c[4], b[8], b[9]);
	or n005(c[5], b[10],b[11]);
	or n006(c[6], b[12],b[13]);
	or n007(c[7], b[14],b[15]);
	
	or n0000(d[0], c[0], c[1]);
	or n0001(d[1], c[3], c[2]);
	or n0002(d[2], c[4], c[5]);
	or n0003(d[3], c[6], c[7]);
	
	or n00000(e[0], d[0], d[1]);
	or n00001(e[1], d[3], d[2]);
	
	or n000000(out, e[0], e[1]);
	
endmodule
