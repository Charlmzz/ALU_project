module not_gate32(a, y);
	output [31:0] a;
	input [31:0] y;
	
	not n0(a[0], y[0]);
	not n1(a[1], y[1]);
	not n2(a[2], y[2]);
	not n3(a[3], y[3]);
	not n4(a[4], y[4]);
	not n5(a[5], y[5]);
	not n6(a[6], y[6]);
	not n7(a[7], y[7]);
	not n8(a[8], y[8]);
	not n9(a[9], y[9]);
	not n10(a[10], y[10]);
	not n11(a[11], y[11]);
	not n12(a[12], y[12]);
	not n13(a[13], y[13]);
	not n14(a[14], y[14]);
	not n15(a[15], y[15]);
	
	not n16(a[16], y[16]);
	not n17(a[17], y[17]);
	not n18(a[18], y[18]);
	not n19(a[19], y[19]);
	not n20(a[20], y[20]);
	not n21(a[21], y[21]);
	not n22(a[22], y[22]);
	not n23(a[23], y[23]);
	not n24(a[24], y[24]);
	not n25(a[25], y[25]);
	not n26(a[26], y[26]);
	not n27(a[27], y[27]);
	not n28(a[28], y[28]);
	not n29(a[29], y[29]);
	not n30(a[30], y[30]);
	not n31(a[31], y[31]);
	
endmodule
